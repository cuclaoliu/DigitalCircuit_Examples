--SHIFT 8BIT 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY SHIFT1 IS 
PORT (
	CLK,RST : IN STD_LOGIC;
	DIN: IN STD_LOGIC;
	QOUT : OUT STD_LOGIC);
END SHIFT1 ;

ARCHITECTURE RTL OF SHIFT1 IS 
SIGNAL REGS : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
  PROCESS (CLK,RST)
  BEGIN
    IF RST='0' THEN REGS<="00000";QOUT<='0';
    ELSIF CLK'EVENT AND CLK='1' THEN 
		REGS(0)<=DIN;
		REGS(1)<=REGS(0);
		REGS(2)<=REGS(1);
		REGS(3)<=REGS(2);
		REGS(4)<=REGS(3);
		QOUT <= REGS(4);
	END IF;
  END PROCESS; 
END RTL;