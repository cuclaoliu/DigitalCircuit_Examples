LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
package mypack is

	subtype BCD is integer range 0 to 9;
	subtype SSD	is STD_LOGIC_VECTOR(0 TO 6);
	
end mypack;
